`default_nettype none
module font (
	xidx,
	yidx,
	char,
	pixel
);
	input wire [3:0] xidx;
	input wire [3:0] yidx;
	input wire [7:0] char;
	output reg pixel;
	always @(*)
		case (char)
			8'd32: pixel = 0;
			8'd33: pixel = ((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd34: pixel = ((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4));
			8'd35: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd36: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 5) && (yidx == 0))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd37: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd38: pixel = (((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd39: pixel = ((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4));
			8'd40: pixel = ((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd41: pixel = ((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd42: pixel = ((((((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd43: pixel = ((((((((((((((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9));
			8'd44: pixel = ((((((((xidx == 3) && (yidx == 8)) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11));
			8'd45: pixel = ((((((((xidx == 0) && (yidx == 6)) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6));
			8'd46: pixel = ((((xidx == 3) && (yidx == 9)) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd47: pixel = ((((((((((((((xidx == 7) && (yidx == 2)) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9));
			8'd48: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd49: pixel = (((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd50: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd51: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd52: pixel = ((((((((((((((((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd53: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd54: pixel = ((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd55: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd56: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd57: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd58: pixel = ((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9));
			8'd59: pixel = ((((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10));
			8'd60: pixel = ((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd61: pixel = ((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd62: pixel = ((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10));
			8'd63: pixel = (((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd64: pixel = (((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd65: pixel = (((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd66: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd67: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd68: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd69: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd70: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd71: pixel = (((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd72: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd73: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd74: pixel = ((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd75: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd76: pixel = ((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd77: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd78: pixel = (((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd79: pixel = ((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd80: pixel = (((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd81: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11));
			8'd82: pixel = ((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd83: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd84: pixel = ((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd85: pixel = (((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd86: pixel = ((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd87: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd88: pixel = ((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd89: pixel = ((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd90: pixel = ((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd91: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd92: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 7) && (yidx == 10));
			8'd93: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd94: pixel = ((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3));
			8'd95: pixel = ((((((((xidx == 0) && (yidx == 12)) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd96: pixel = ((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2));
			8'd97: pixel = ((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd98: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd99: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd100: pixel = ((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd101: pixel = (((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd102: pixel = (((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd103: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd104: pixel = (((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd105: pixel = (((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd106: pixel = (((((((((((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd107: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd108: pixel = (((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd109: pixel = (((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd110: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd111: pixel = ((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd112: pixel = ((((((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12));
			8'd113: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd114: pixel = ((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd115: pixel = ((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd116: pixel = ((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd117: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd118: pixel = ((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd119: pixel = ((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd120: pixel = ((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd121: pixel = ((((((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd122: pixel = ((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd123: pixel = (((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd124: pixel = ((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd125: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10));
			8'd126: pixel = ((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3));
			default: pixel = 0;
		endcase
endmodule
module font_cp437 (
	xidx,
	yidx,
	char,
	pixel
);
	input wire [3:0] xidx;
	input wire [3:0] yidx;
	input wire [7:0] char;
	output reg pixel;
	always @(*)
		case (char)
			8'd0: pixel = 0;
			8'd1: pixel = ((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd2: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd3: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 3)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 4) && (yidx == 10));
			8'd4: pixel = (((((((((((((((((((((((((xidx == 4) && (yidx == 3)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9));
			8'd5: pixel = ((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd6: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd7: pixel = ((((((((((((xidx == 3) && (yidx == 5)) || ((xidx == 4) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8));
			8'd8: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 2) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13));
			8'd9: pixel = ((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9));
			8'd10: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 2) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13));
			8'd11: pixel = (((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd12: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd13: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10));
			8'd14: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11));
			8'd15: pixel = ((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd16: pixel = (((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 1) && (yidx == 10));
			8'd17: pixel = (((((((((((((((((((((((((((((xidx == 7) && (yidx == 2)) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 7) && (yidx == 10));
			8'd18: pixel = ((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd19: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd20: pixel = (((((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd21: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12));
			8'd22: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 8)) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd23: pixel = ((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11));
			8'd24: pixel = ((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd25: pixel = ((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd26: pixel = (((((((((((((((xidx == 4) && (yidx == 4)) || ((xidx == 5) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8));
			8'd27: pixel = (((((((((((((((xidx == 3) && (yidx == 4)) || ((xidx == 4) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8));
			8'd28: pixel = (((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8));
			8'd29: pixel = ((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8));
			8'd30: pixel = (((((((((((((((((((((((((((((((xidx == 4) && (yidx == 3)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9));
			8'd31: pixel = (((((((((((((((((((((((((((((((xidx == 1) && (yidx == 3)) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9));
			8'd32: pixel = 0;
			8'd33: pixel = ((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd34: pixel = ((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4));
			8'd35: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd36: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 5) && (yidx == 0))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd37: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd38: pixel = (((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd39: pixel = ((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4));
			8'd40: pixel = ((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd41: pixel = ((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd42: pixel = ((((((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd43: pixel = ((((((((((((((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9));
			8'd44: pixel = ((((((((xidx == 3) && (yidx == 8)) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11));
			8'd45: pixel = ((((((((xidx == 0) && (yidx == 6)) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6));
			8'd46: pixel = ((((xidx == 3) && (yidx == 9)) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd47: pixel = ((((((((((((((xidx == 7) && (yidx == 2)) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9));
			8'd48: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd49: pixel = (((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd50: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd51: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd52: pixel = ((((((((((((((((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd53: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd54: pixel = ((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd55: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd56: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd57: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd58: pixel = ((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9));
			8'd59: pixel = ((((((((((xidx == 3) && (yidx == 3)) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10));
			8'd60: pixel = ((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd61: pixel = ((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd62: pixel = ((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10));
			8'd63: pixel = (((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd64: pixel = (((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd65: pixel = (((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd66: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd67: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd68: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd69: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd70: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd71: pixel = (((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd72: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd73: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd74: pixel = ((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd75: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd76: pixel = ((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd77: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd78: pixel = (((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd79: pixel = ((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd80: pixel = (((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd81: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11));
			8'd82: pixel = ((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd83: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd84: pixel = ((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd85: pixel = (((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd86: pixel = ((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd87: pixel = ((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd88: pixel = ((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd89: pixel = ((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd90: pixel = ((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd91: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd92: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 7) && (yidx == 10));
			8'd93: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd94: pixel = ((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3));
			8'd95: pixel = ((((((((xidx == 0) && (yidx == 12)) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd96: pixel = ((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2));
			8'd97: pixel = ((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd98: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd99: pixel = ((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd100: pixel = ((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd101: pixel = (((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd102: pixel = (((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd103: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd104: pixel = (((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd105: pixel = (((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd106: pixel = (((((((((((((((((((((((((((xidx == 5) && (yidx == 2)) || ((xidx == 6) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd107: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd108: pixel = (((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd109: pixel = (((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd110: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd111: pixel = ((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd112: pixel = ((((((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12));
			8'd113: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd114: pixel = ((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd115: pixel = ((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd116: pixel = ((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd117: pixel = (((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd118: pixel = ((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd119: pixel = ((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd120: pixel = ((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd121: pixel = ((((((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd122: pixel = ((((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd123: pixel = (((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd124: pixel = ((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd125: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10));
			8'd126: pixel = ((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3));
			8'd127: pixel = (((((((((((((((((((((((xidx == 4) && (yidx == 4)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9));
			8'd128: pixel = (((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12));
			8'd129: pixel = (((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd130: pixel = (((((((((((((((((((((((((((((((((xidx == 5) && (yidx == 1)) || ((xidx == 6) && (yidx == 1))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd131: pixel = ((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd132: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd133: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd134: pixel = ((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 1)) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd135: pixel = ((((((((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11));
			8'd136: pixel = (((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd137: pixel = (((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd138: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd139: pixel = (((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd140: pixel = (((((((((((((((((((((((((xidx == 3) && (yidx == 1)) || ((xidx == 4) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd141: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd142: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd143: pixel = ((((((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd144: pixel = (((((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 5) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd145: pixel = (((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd146: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd147: pixel = ((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd148: pixel = ((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd149: pixel = ((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd150: pixel = (((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 1)) || ((xidx == 4) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd151: pixel = (((((((((((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd152: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12));
			8'd153: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd154: pixel = (((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd155: pixel = ((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 1)) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd156: pixel = (((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 1)) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd157: pixel = ((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 2)) || ((xidx == 1) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd158: pixel = ((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 1)) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd159: pixel = ((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12));
			8'd160: pixel = ((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd161: pixel = (((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd162: pixel = ((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd163: pixel = (((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd164: pixel = (((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd165: pixel = (((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd166: pixel = (((((((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6));
			8'd167: pixel = (((((((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6));
			8'd168: pixel = (((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd169: pixel = (((((((((((((xidx == 1) && (yidx == 6)) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9));
			8'd170: pixel = (((((((((((((xidx == 1) && (yidx == 6)) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9));
			8'd171: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd172: pixel = (((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12));
			8'd173: pixel = ((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd174: pixel = ((((((((((((((((((((xidx == 3) && (yidx == 4)) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8));
			8'd175: pixel = ((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8));
			8'd176: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 7) && (yidx == 0))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 5) && (yidx == 13));
			8'd177: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd178: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13));
			8'd179: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd180: pixel = (((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd181: pixel = ((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd182: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd183: pixel = (((((((((((((((((((((((((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd184: pixel = ((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd185: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd186: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd187: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd188: pixel = (((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7));
			8'd189: pixel = (((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7));
			8'd190: pixel = ((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7));
			8'd191: pixel = (((((((((((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd192: pixel = ((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd193: pixel = (((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd194: pixel = (((((((((((((((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd195: pixel = ((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd196: pixel = (((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd197: pixel = (((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd198: pixel = ((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd199: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd200: pixel = (((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd201: pixel = (((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd202: pixel = (((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd203: pixel = (((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd204: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd205: pixel = ((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd206: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd207: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd208: pixel = (((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd209: pixel = ((((((((((((((((((((((((((((((xidx == 0) && (yidx == 5)) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd210: pixel = (((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd211: pixel = (((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd212: pixel = ((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7));
			8'd213: pixel = ((((((((((((((((((((((((((xidx == 3) && (yidx == 5)) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd214: pixel = (((((((((((((((((((((((((((((((xidx == 2) && (yidx == 7)) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd215: pixel = (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 0)) || ((xidx == 3) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13));
			8'd216: pixel = ((((((((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd217: pixel = (((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7));
			8'd218: pixel = ((((((((((((((((((xidx == 3) && (yidx == 7)) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd219: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 2) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 8) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 8) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 8) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 8) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 8) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 8) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 8) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 8) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 8) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 8) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 8) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13))) || ((xidx == 8) && (yidx == 13));
			8'd220: pixel = (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 7)) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 8) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 8) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 8) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 8) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 8) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13))) || ((xidx == 8) && (yidx == 13));
			8'd221: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 2) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 0) && (yidx == 11))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 0) && (yidx == 12))) || ((xidx == 1) && (yidx == 12))) || ((xidx == 2) && (yidx == 12))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 0) && (yidx == 13))) || ((xidx == 1) && (yidx == 13))) || ((xidx == 2) && (yidx == 13))) || ((xidx == 3) && (yidx == 13));
			8'd222: pixel = ((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 4) && (yidx == 0)) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 8) && (yidx == 0))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 8) && (yidx == 1))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 8) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 8) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 8) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 8) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 8) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 8) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 8) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10))) || ((xidx == 8) && (yidx == 10))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 5) && (yidx == 11))) || ((xidx == 6) && (yidx == 11))) || ((xidx == 7) && (yidx == 11))) || ((xidx == 8) && (yidx == 11))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 5) && (yidx == 12))) || ((xidx == 6) && (yidx == 12))) || ((xidx == 7) && (yidx == 12))) || ((xidx == 8) && (yidx == 12))) || ((xidx == 4) && (yidx == 13))) || ((xidx == 5) && (yidx == 13))) || ((xidx == 6) && (yidx == 13))) || ((xidx == 7) && (yidx == 13))) || ((xidx == 8) && (yidx == 13));
			8'd223: pixel = (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((xidx == 0) && (yidx == 0)) || ((xidx == 1) && (yidx == 0))) || ((xidx == 2) && (yidx == 0))) || ((xidx == 3) && (yidx == 0))) || ((xidx == 4) && (yidx == 0))) || ((xidx == 5) && (yidx == 0))) || ((xidx == 6) && (yidx == 0))) || ((xidx == 7) && (yidx == 0))) || ((xidx == 8) && (yidx == 0))) || ((xidx == 0) && (yidx == 1))) || ((xidx == 1) && (yidx == 1))) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 8) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 8) && (yidx == 2))) || ((xidx == 0) && (yidx == 3))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 8) && (yidx == 3))) || ((xidx == 0) && (yidx == 4))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 8) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 8) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 8) && (yidx == 6));
			8'd224: pixel = ((((((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd225: pixel = ((((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11))) || ((xidx == 2) && (yidx == 12));
			8'd226: pixel = (((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10));
			8'd227: pixel = (((((((((((((((((((((((((((((((xidx == 1) && (yidx == 4)) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd228: pixel = ((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 7) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd229: pixel = (((((((((((((((((((((((((xidx == 2) && (yidx == 5)) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd230: pixel = (((((((((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 1) && (yidx == 11))) || ((xidx == 2) && (yidx == 11));
			8'd231: pixel = ((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd232: pixel = ((((((((((((((((((((((((((((((((((((xidx == 1) && (yidx == 2)) || ((xidx == 2) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd233: pixel = (((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd234: pixel = (((((((((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd235: pixel = (((((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd236: pixel = ((((((((((((((((((((((((xidx == 1) && (yidx == 5)) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd237: pixel = ((((((((((((((((((((((((((((((((((((((xidx == 6) && (yidx == 2)) || ((xidx == 7) && (yidx == 2))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10));
			8'd238: pixel = (((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd239: pixel = (((((((((((((((((((((((((((((((((xidx == 2) && (yidx == 3)) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 7) && (yidx == 8))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd240: pixel = (((((((((((((((((((((xidx == 1) && (yidx == 3)) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9))) || ((xidx == 7) && (yidx == 9));
			8'd241: pixel = ((((((((((((((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 7) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 0) && (yidx == 10))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10))) || ((xidx == 7) && (yidx == 10));
			8'd242: pixel = ((((((((((((((((((((xidx == 2) && (yidx == 2)) || ((xidx == 3) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd243: pixel = ((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10))) || ((xidx == 6) && (yidx == 10));
			8'd244: pixel = (((((((((((((((((((((((((((((xidx == 4) && (yidx == 2)) || ((xidx == 5) && (yidx == 2))) || ((xidx == 6) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 6) && (yidx == 3))) || ((xidx == 7) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 3) && (yidx == 11))) || ((xidx == 4) && (yidx == 11))) || ((xidx == 3) && (yidx == 12))) || ((xidx == 4) && (yidx == 12))) || ((xidx == 3) && (yidx == 13))) || ((xidx == 4) && (yidx == 13));
			8'd245: pixel = (((((((((((((((((((((((((((xidx == 3) && (yidx == 0)) || ((xidx == 4) && (yidx == 0))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 0) && (yidx == 8))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 0) && (yidx == 9))) || ((xidx == 1) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 1) && (yidx == 10))) || ((xidx == 2) && (yidx == 10))) || ((xidx == 3) && (yidx == 10));
			8'd246: pixel = ((((((((((((((((xidx == 3) && (yidx == 2)) || ((xidx == 4) && (yidx == 2))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 7) && (yidx == 6))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10));
			8'd247: pixel = ((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 7) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 7) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8));
			8'd248: pixel = ((((((((((((((xidx == 2) && (yidx == 1)) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4));
			8'd249: pixel = ((((xidx == 3) && (yidx == 6)) || ((xidx == 4) && (yidx == 6))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7));
			8'd250: pixel = ((xidx == 3) && (yidx == 7)) || ((xidx == 4) && (yidx == 7));
			8'd251: pixel = ((((((((((((((((((((((((((((((xidx == 4) && (yidx == 1)) || ((xidx == 5) && (yidx == 1))) || ((xidx == 6) && (yidx == 1))) || ((xidx == 7) && (yidx == 1))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 0) && (yidx == 7))) || ((xidx == 1) && (yidx == 7))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 1) && (yidx == 8))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 3) && (yidx == 10))) || ((xidx == 4) && (yidx == 10))) || ((xidx == 5) && (yidx == 10));
			8'd252: pixel = ((((((((((((((((((((((((xidx == 0) && (yidx == 1)) || ((xidx == 1) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 4) && (yidx == 1))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 2) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 5) && (yidx == 2))) || ((xidx == 1) && (yidx == 3))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 4) && (yidx == 3))) || ((xidx == 5) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6));
			8'd253: pixel = (((((((((((((((((((xidx == 1) && (yidx == 1)) || ((xidx == 2) && (yidx == 1))) || ((xidx == 3) && (yidx == 1))) || ((xidx == 0) && (yidx == 2))) || ((xidx == 1) && (yidx == 2))) || ((xidx == 3) && (yidx == 2))) || ((xidx == 4) && (yidx == 2))) || ((xidx == 2) && (yidx == 3))) || ((xidx == 3) && (yidx == 3))) || ((xidx == 1) && (yidx == 4))) || ((xidx == 2) && (yidx == 4))) || ((xidx == 0) && (yidx == 5))) || ((xidx == 1) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 0) && (yidx == 6))) || ((xidx == 1) && (yidx == 6))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6));
			8'd254: pixel = ((((((((((((((((((((((((((((((xidx == 2) && (yidx == 4)) || ((xidx == 3) && (yidx == 4))) || ((xidx == 4) && (yidx == 4))) || ((xidx == 5) && (yidx == 4))) || ((xidx == 6) && (yidx == 4))) || ((xidx == 2) && (yidx == 5))) || ((xidx == 3) && (yidx == 5))) || ((xidx == 4) && (yidx == 5))) || ((xidx == 5) && (yidx == 5))) || ((xidx == 6) && (yidx == 5))) || ((xidx == 2) && (yidx == 6))) || ((xidx == 3) && (yidx == 6))) || ((xidx == 4) && (yidx == 6))) || ((xidx == 5) && (yidx == 6))) || ((xidx == 6) && (yidx == 6))) || ((xidx == 2) && (yidx == 7))) || ((xidx == 3) && (yidx == 7))) || ((xidx == 4) && (yidx == 7))) || ((xidx == 5) && (yidx == 7))) || ((xidx == 6) && (yidx == 7))) || ((xidx == 2) && (yidx == 8))) || ((xidx == 3) && (yidx == 8))) || ((xidx == 4) && (yidx == 8))) || ((xidx == 5) && (yidx == 8))) || ((xidx == 6) && (yidx == 8))) || ((xidx == 2) && (yidx == 9))) || ((xidx == 3) && (yidx == 9))) || ((xidx == 4) && (yidx == 9))) || ((xidx == 5) && (yidx == 9))) || ((xidx == 6) && (yidx == 9));
			8'd255: pixel = 0;
			default: pixel = 0;
		endcase
endmodule
module sim;
	reg clock;
	wire MDA_HSYNC;
	wire MDA_VSYNC;
	wire MDA_DATA;
	wire MDA_INTENSITY;
	mda_core dut(
		.clock(clock),
		.MDA_HSYNC(MDA_HSYNC),
		.MDA_VSYNC(MDA_VSYNC),
		.MDA_DATA(MDA_DATA),
		.MDA_INTENSITY(MDA_INTENSITY)
	);
	initial begin
		clock = 0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < 600000; i = i + 1)
				begin
					clock = !clock;
					#(5)
						;
					clock = !clock;
					#(5)
						;
				end
		end
		$dumpvars(1, sim);
		$dumpfile("out.vcd");
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < 900000; i = i + 1)
				begin
					clock = !clock;
					#(5)
						;
					clock = !clock;
					#(5)
						;
				end
		end
	end
endmodule
module mda_core (
	clock,
	MDA_HSYNC,
	MDA_VSYNC,
	MDA_DATA,
	MDA_INTENSITY
);
	input wire clock;
	output wire MDA_HSYNC;
	output wire MDA_VSYNC;
	output wire MDA_DATA;
	output wire MDA_INTENSITY;
	reg mda_hsync_int = 'h0;
	reg mda_vsync_int = 'h0;
	reg mda_intensity_int = 'h0;
	reg mda_shifter_load = 'h0;
	reg [30:0] ctr;
	reg inv;
	reg [8:0] yctr = 'h0;
	reg [15:0] xctr = 'h0;
	assign MDA_HSYNC = mda_hsync_int;
	assign MDA_VSYNC = mda_vsync_int;
	wire valid = ((xctr >= 17) && (xctr < 737)) && (yctr < 350);
	wire m_bit;
	reg [6:0] xchar;
	reg [6:0] ychar;
	reg [6:0] xchar_ctr;
	reg [6:0] ychar_ctr;
	reg [7:0] char;
	always @(*) begin
		char = 0;
		if ((xchar < 64) && (ychar < 4))
			char = {ychar[1:0], xchar[5:0]};
	end
	font_cp437 thefont(
		.xidx(xchar_ctr),
		.yidx(ychar_ctr),
		.char(char),
		.pixel(m_bit)
	);
	assign MDA_DATA = m_bit && valid;
	assign MDA_INTENSITY = valid;
	always @(posedge clock) begin
		ctr <= ctr + 1;
		if ((ctr >= 48000000) && (mda_vsync_int == 0)) begin
			ctr <= 0;
			inv <= !inv;
		end
		xchar_ctr <= xchar_ctr + 1;
		if (xchar_ctr == 8) begin
			xchar_ctr <= 0;
			xchar <= xchar + 1;
		end
		if (!valid) begin
			xchar_ctr <= 0;
			xchar <= 0;
		end
		xctr <= xctr + 1'b1;
		case (xctr)
			'd748: mda_hsync_int <= 1'b1;
			'd883: begin
				mda_hsync_int <= 1'b0;
				yctr <= yctr + 1'b1;
				ychar_ctr <= ychar_ctr + 1;
				if (ychar_ctr == 13) begin
					ychar_ctr <= 0;
					ychar <= ychar + 1;
				end
				xctr <= 'd0;
				if (yctr == 'd348)
					mda_vsync_int <= 1'b0;
				if (yctr == 'd364)
					mda_vsync_int <= 1'b1;
				if (yctr == 'd368) begin
					yctr <= 'h0;
					ychar <= 0;
					ychar_ctr <= 0;
				end
			end
			default:
				;
		endcase
	end
endmodule
